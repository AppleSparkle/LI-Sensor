// Copyright (C) 1991-2012 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 12.1 Build 177 11/07/2012 SJ Full Version
// Created on Fri Jun 21 15:48:10 2013

// synthesis message_off 10175

`timescale 1ns/1ns

module syst_ctrl_statemachine (
    reset,clock,C1,C2,C3,C4,C5,C6,C7,C8,C9,C10,C11,C12,START,
    C1_EN,C2_EN,C3_EN,C4_EN,C5_EN,C6_EN,C7_EN,C8_EN,C9_EN,C10_EN,C11_EN,C12_EN,CLR);

    input reset;
    input clock;
    input C1;
    input C2;
    input C3;
    input C4;
    input C5;
    input C6;
    input C7;
    input C8;
    input C9;
    input C10;
    input C11;
    input C12;
    input START;
    tri0 reset;
    tri0 C1;
    tri0 C2;
    tri0 C3;
    tri0 C4;
    tri0 C5;
    tri0 C6;
    tri0 C7;
    tri0 C8;
    tri0 C9;
    tri0 C10;
    tri0 C11;
    tri0 C12;
    tri0 START;
    output C1_EN;
    output C2_EN;
    output C3_EN;
    output C4_EN;
    output C5_EN;
    output C6_EN;
    output C7_EN;
    output C8_EN;
    output C9_EN;
    output C10_EN;
    output C11_EN;
    output C12_EN;
    output CLR;
    reg C1_EN;
    reg reg_C1_EN;
    reg C2_EN;
    reg reg_C2_EN;
    reg C3_EN;
    reg reg_C3_EN;
    reg C4_EN;
    reg reg_C4_EN;
    reg C5_EN;
    reg reg_C5_EN;
    reg C6_EN;
    reg reg_C6_EN;
    reg C7_EN;
    reg reg_C7_EN;
    reg C8_EN;
    reg reg_C8_EN;
    reg C9_EN;
    reg reg_C9_EN;
    reg C10_EN;
    reg reg_C10_EN;
    reg C11_EN;
    reg reg_C11_EN;
    reg C12_EN;
    reg reg_C12_EN;
    reg CLR;
    reg reg_CLR;
    reg [13:0] fstate;
    reg [13:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3,state5=4,state6=5,state7=6,state8=7,state9=8,state10=9,state11=10,state12=11,state13=12,state14=13;

    initial
    begin
        reg_C1_EN <= 1'b0;
        reg_C2_EN <= 1'b0;
        reg_C3_EN <= 1'b0;
        reg_C4_EN <= 1'b0;
        reg_C5_EN <= 1'b0;
        reg_C6_EN <= 1'b0;
        reg_C7_EN <= 1'b0;
        reg_C8_EN <= 1'b0;
        reg_C9_EN <= 1'b0;
        reg_C10_EN <= 1'b0;
        reg_C11_EN <= 1'b0;
        reg_C12_EN <= 1'b0;
        reg_CLR <= 1'b0;
    end

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
            C1_EN <= reg_C1_EN;
            C2_EN <= reg_C2_EN;
            C3_EN <= reg_C3_EN;
            C4_EN <= reg_C4_EN;
            C5_EN <= reg_C5_EN;
            C6_EN <= reg_C6_EN;
            C7_EN <= reg_C7_EN;
            C8_EN <= reg_C8_EN;
            C9_EN <= reg_C9_EN;
            C10_EN <= reg_C10_EN;
            C11_EN <= reg_C11_EN;
            C12_EN <= reg_C12_EN;
            CLR <= reg_CLR;
        end
    end

    always @(fstate or reset or C1 or C2 or C3 or C4 or C5 or C6 or C7 or C8 or C9 or C10 or C11 or C12 or START)
    begin
        if (reset) begin
            reg_fstate <= state1;
            reg_C1_EN <= 1'b0;
            reg_C2_EN <= 1'b0;
            reg_C3_EN <= 1'b0;
            reg_C4_EN <= 1'b0;
            reg_C5_EN <= 1'b0;
            reg_C6_EN <= 1'b0;
            reg_C7_EN <= 1'b0;
            reg_C8_EN <= 1'b0;
            reg_C9_EN <= 1'b0;
            reg_C10_EN <= 1'b0;
            reg_C11_EN <= 1'b0;
            reg_C12_EN <= 1'b0;
            reg_CLR <= 1'b0;
        end
        else begin
            reg_C1_EN <= 1'b0;
            reg_C2_EN <= 1'b0;
            reg_C3_EN <= 1'b0;
            reg_C4_EN <= 1'b0;
            reg_C5_EN <= 1'b0;
            reg_C6_EN <= 1'b0;
            reg_C7_EN <= 1'b0;
            reg_C8_EN <= 1'b0;
            reg_C9_EN <= 1'b0;
            reg_C10_EN <= 1'b0;
            reg_C11_EN <= 1'b0;
            reg_C12_EN <= 1'b0;
            reg_CLR <= 1'b0;
            case (fstate)
                state1: begin
                    if (~(START))
                        reg_fstate <= state1;
                    else if (START)
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;
                end
                state2: begin
                    if (~(C1))
                        reg_fstate <= state2;
                    else if (C1)
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    reg_C1_EN <= 1'b1;
                end
                state3: begin
                    if (~(C2))
                        reg_fstate <= state3;
                    else if (C2)
                        reg_fstate <= state4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    reg_C2_EN <= 1'b1;
                end
                state4: begin
                    if (~(C3))
                        reg_fstate <= state4;
                    else if (C3)
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    reg_C3_EN <= 1'b1;
                end
                state5: begin
                    if (~(C4))
                        reg_fstate <= state5;
                    else if (C4)
                        reg_fstate <= state6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    reg_C4_EN <= 1'b1;
                end
                state6: begin
                    if (~(C5))
                        reg_fstate <= state6;
                    else if (C5)
                        reg_fstate <= state7;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state6;

                    reg_C5_EN <= 1'b1;
                end
                state7: begin
                    if (~(C6))
                        reg_fstate <= state7;
                    else if (C6)
                        reg_fstate <= state8;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state7;

                    reg_C6_EN <= 1'b1;
                end
                state8: begin
                    if (~(C7))
                        reg_fstate <= state8;
                    else if (C7)
                        reg_fstate <= state9;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state8;

                    reg_C7_EN <= 1'b1;
                end
                state9: begin
                    if (~(C8))
                        reg_fstate <= state9;
                    else if (C8)
                        reg_fstate <= state10;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state9;

                    reg_C8_EN <= 1'b1;
                end
                state10: begin
                    if (C9)
                        reg_fstate <= state11;
                    else if (~(C9))
                        reg_fstate <= state10;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state10;

                    reg_C9_EN <= 1'b1;
                end
                state11: begin
                    if (C10)
                        reg_fstate <= state12;
                    else if (~(C10))
                        reg_fstate <= state11;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state11;

                    reg_C10_EN <= 1'b1;
                end
                state12: begin
                    if (~(C11))
                        reg_fstate <= state12;
                    else if (C11)
                        reg_fstate <= state13;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state12;

                    reg_C11_EN <= 1'b1;
                end
                state13: begin
                    if (~(C12))
                        reg_fstate <= state13;
                    else if (C12)
                        reg_fstate <= state14;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state13;

                    reg_C12_EN <= 1'b1;
                end
                state14: begin
                    reg_fstate <= state1;

                    reg_CLR <= 1'b1;
                end
                default: begin
                    reg_C1_EN <= 1'bx;
                    reg_C2_EN <= 1'bx;
                    reg_C3_EN <= 1'bx;
                    reg_C4_EN <= 1'bx;
                    reg_C5_EN <= 1'bx;
                    reg_C6_EN <= 1'bx;
                    reg_C7_EN <= 1'bx;
                    reg_C8_EN <= 1'bx;
                    reg_C9_EN <= 1'bx;
                    reg_C10_EN <= 1'bx;
                    reg_C11_EN <= 1'bx;
                    reg_C12_EN <= 1'bx;
                    reg_CLR <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // syst_ctrl_statemachine
